module main;
    initial $hello;
endmodule